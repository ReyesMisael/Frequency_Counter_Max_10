library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Empty_Buf is 

port (
		Z : in std_logic_vector(7 to 0) 
		);

end entity;

architecture Arch of Empty_buf is
	begin
	

end Arch;